module InstrMem (input [31:0]address, output [31:0]data,output [5:0]lookahead);
  reg [7:0] mem [0:63];
  wire [7:0]w;
  initial begin
    mem[0]=8'b 00000000;
    mem[1]=8'b 00100010;
    mem[2]=8'b 00100000;
    mem[3]=8'b 00000001;
    mem[4]=8'b 00001100;
    mem[5]=8'b 00000000;
    mem[6]=8'b 00000000;
    mem[7]=8'b 00000000;
    mem[8]=8'b 00000000;
    mem[9]=8'b 00100010;
    mem[10]=8'b 00101000;
    mem[11]=8'b 00000000;
    mem[12]=8'b 00000000;
    mem[13]=8'b 00100010;
    mem[14]=8'b 00110000;
    mem[15]=8'b 00000010;
    mem[16]=8'b 00000000; //rtype
    mem[17]=8'b 00100010;
    mem[18]=8'b 00111000;
    mem[19]=8'b 00000001;
    //mem[20]=8'b 00001100; //Exm
    //mem[21]=8'b 00000000;
    //mem[22]=8'b 00000000;
    //mem[23]=8'b 00000000;
    //mem[20]=8'b 00000100; //jump 28
    //mem[21]=8'b 00000000;
    //mem[22]=8'b 00000000;
    //mem[23]=8'b 00000111;
    mem[20]=8'b 00000000; //rtype
    mem[21]=8'b 00100011;
    mem[22]=8'b 01000000;
    mem[23]=8'b 00000000;
    mem[24]=8'b 00000000; //rtype
    mem[25]=8'b 00100011;
    mem[26]=8'b 01000000;
    mem[27]=8'b 00000000;
    mem[28]=8'b 00010000; //Exr
    mem[29]=8'b 01100100;
    mem[30]=8'b 01001000;
    mem[31]=8'b 00000000;
    //mem[28]=8'b 00000000; //rtype
    //mem[29]=8'b 01000001;
    //mem[30]=8'b 00011000;
    //mem[31]=8'b 00000000;
    mem[32]=8'b 00000000; //rtype
    mem[33]=8'b 00000001;
    mem[34]=8'b 00000010;
    mem[35]=8'b 00000011;
    //mem[36]=8'b 00001010; //jr
    //mem[37]=8'b 00000001;
    //mem[38]=8'b 00000110;
    //mem[39]=8'b 00000111;
    mem[36]=8'b 00000000; //rtype
    mem[37]=8'b 00000001;
    mem[38]=8'b 00000010;
    mem[39]=8'b 00000011;
    mem[40]=8'b 00000000; //rtype
    mem[41]=8'b 00000001;
    mem[42]=8'b 00000010;
    mem[43]=8'b 00000011;
    mem[44]=8'b 00000000; //rtype
    mem[45]=8'b 00000101;
    mem[46]=8'b 00000110;
    mem[47]=8'b 00000111;
    mem[48]=8'b 00000000;
    mem[49]=8'b 00000001;
    mem[50]=8'b 00000010;
    mem[51]=8'b 00000011;
    mem[52]=8'b 00000100;
    mem[53]=8'b 00000101;
    mem[54]=8'b 00000110;
    mem[55]=8'b 00000111;
    mem[56]=8'b 00000000;
    mem[57]=8'b 00000001;
    mem[58]=8'b 00000010;
    mem[59]=8'b 00000011;
    mem[60]=8'b 00000100;
    mem[61]=8'b 00000101;
    mem[62]=8'b 00000110;
    mem[63]=8'b 00000111;
end
wire [31:0]address1,address2,address3;
CSA_32bit f1 (address,32'b00000000000000000000000000000001,1'b0,address1,co,ov),
          f2 (address,32'b00000000000000000000000000000010,1'b0,address2,co,ov),
          f3 (address,32'b00000000000000000000000000000011,1'b0,address3,co,ov);
assign data[31:24]=mem[address];
assign data[23:16]=mem[address1];
assign data[15:8]=mem[address2];
assign data[7:0]=mem[address3];
assign w=mem[address+4];
assign lookahead=w[7:2];
endmodule