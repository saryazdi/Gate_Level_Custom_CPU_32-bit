module RegisterFile (input [4:0]ReadAd1,ReadAd2,WRdst,input [31:0]WRdata0, input wr,wr1,clk, output [31:0]ReadData1,ReadData2,ReadData3);
wire [4:0] Wr1Ad1;
wire [31:0]en,Exr,EN,EN1;
wire [31:0]s31,s30,s29,s28,s27,s26,s25,s24,s23,s22,s21,s20,s19,s18,s17,s16,s15,s14,s13,s12,s11,s10,s9,s8,s7,s6,s5,s4,s3,s2,s1,s0,c;
wire [31:0]WrData31,WrData30,WrData29,WrData28,WrData27,WrData26,WrData25,WrData24,WrData23,WrData22,WrData21,WrData20,WrData19,WrData18,WrData17,WrData16,WrData15,WrData14,WrData13,WrData12,WrData11,WrData10,WrData9,WrData8,WrData7,WrData6,WrData5,WrData4,WrData3,WrData2,WrData1;
assign Wr1Ad1 = (wr1) ? ReadAd1 : 5'b00000;
decoder_32bit D0 (WRdst,EN),
              D1 (Wr1Ad1,Exr);
assign EN1=Exr|EN;
assign en=(Exr==32'b00000000000000000000000000000001)? EN: EN1;
reg_32bit R0 (32'b00000000000000000000000000000000,1'b1,1'b1,clk,s0),
          R1 (32'b00000000000000000000000000000101,1'b1,1'b1,clk,s1),
          R2 (32'b00000000000000000000000000000100,1'b1,1'b1,clk,s2),
          R3 (WrData3,en[3],wr,clk,s3),
          R4 (WrData4,en[4],wr,clk,s4),
          R5 (WrData5,en[5],wr,clk,s5),
          R6 (WrData6,en[6],wr,clk,s6),
          R7 (WrData7,en[7],wr,clk,s7),
          R8 (WrData8,en[8],wr,clk,s8),
          R9 (WrData9,en[9],wr,clk,s9),
          R10 (WrData10,en[10],wr,clk,s10),
          R11 (WrData11,en[11],wr,clk,s11),
          R12 (WrData12,en[12],wr,clk,s12),
          R13 (WrData13,en[13],wr,clk,s13),
          R14 (WrData14,en[14],wr,clk,s14),
          R15 (WrData15,en[15],wr,clk,s15),
          R16 (WrData16,en[16],wr,clk,s16),
          R17 (WrData17,en[17],wr,clk,s17),
          R18 (WrData18,en[18],wr,clk,s18),
          R19 (WrData19,en[19],wr,clk,s19),
          R20 (WrData20,en[20],wr,clk,s20),
          R21 (WrData21,en[21],wr,clk,s21),
          R22 (WrData22,en[22],wr,clk,s22),
          R23 (WrData23,en[23],wr,clk,s23),
          R24 (WrData24,en[24],wr,clk,s24),
          R25 (WrData25,en[25],wr,clk,s25),
          R26 (WrData26,en[26],wr,clk,s26),
          R27 (WrData27,en[27],wr,clk,s27),
          R28 (WrData28,en[28],wr,clk,s28),
          R29 (WrData29,en[29],wr,clk,s29),
          R30 (WrData30,en[30],wr,clk,s30),
          R31 (WrData31,en[31],wr,clk,s31);
mux_2x32 o1 (WRdata0,ReadData2,Exr[1],WrData1),
         o2 (WRdata0,ReadData2,Exr[2],WrData2),
         o3 (WRdata0,ReadData2,Exr[3],WrData3),
         o4 (WRdata0,ReadData2,Exr[4],WrData4),
         o5 (WRdata0,ReadData2,Exr[5],WrData5),
         o6 (WRdata0,ReadData2,Exr[6],WrData6),
         o7 (WRdata0,ReadData2,Exr[7],WrData7),
         o8 (WRdata0,ReadData2,Exr[8],WrData8),
         o9 (WRdata0,ReadData2,Exr[9],WrData9),
         o10 (WRdata0,ReadData2,Exr[10],WrData10),
         o11 (WRdata0,ReadData2,Exr[11],WrData11),
         o12 (WRdata0,ReadData2,Exr[12],WrData12),
         o13 (WRdata0,ReadData2,Exr[13],WrData13),
         o14 (WRdata0,ReadData2,Exr[14],WrData14),
         o15 (WRdata0,ReadData2,Exr[15],WrData15),
         o16 (WRdata0,ReadData2,Exr[16],WrData16),
         o17 (WRdata0,ReadData2,Exr[17],WrData17),
         o18 (WRdata0,ReadData2,Exr[18],WrData18),
         o19 (WRdata0,ReadData2,Exr[19],WrData19),
         o20 (WRdata0,ReadData2,Exr[20],WrData20),
         o21 (WRdata0,ReadData2,Exr[21],WrData21),
         o22 (WRdata0,ReadData2,Exr[22],WrData22),
         o23 (WRdata0,ReadData2,Exr[23],WrData23),
         o24 (WRdata0,ReadData2,Exr[24],WrData24),
         o25 (WRdata0,ReadData2,Exr[25],WrData25),
         o26 (WRdata0,ReadData2,Exr[26],WrData26),
         o27 (WRdata0,ReadData2,Exr[27],WrData27),
         o28 (WRdata0,ReadData2,Exr[28],WrData28),
         o29 (WRdata0,ReadData2,Exr[29],WrData29),
         o30 (WRdata0,ReadData2,Exr[30],WrData30),
         o31 (WRdata0,ReadData2,Exr[31],WrData31);
mux_32x1 m0 (s31[0],s30[0],s29[0],s28[0],s27[0],s26[0],s25[0],s24[0],s23[0],s22[0],s21[0],s20[0],s19[0],s18[0],s17[0],s16[0],s15[0],s14[0],s13[0],s12[0],s11[0],s10[0],s9[0],s8[0],s7[0],s6[0],s5[0],s4[0],s3[0],s2[0],s1[0],s0[0],ReadAd1,ReadData1[0]),
         m1 (s31[1],s30[1],s29[1],s28[1],s27[1],s26[1],s25[1],s24[1],s23[1],s22[1],s21[1],s20[1],s19[1],s18[1],s17[1],s16[1],s15[1],s14[1],s13[1],s12[1],s11[1],s10[1],s9[1],s8[1],s7[1],s6[1],s5[1],s4[1],s3[1],s2[1],s1[1],s0[1],ReadAd1,ReadData1[1]),
         m2 (s31[2],s30[2],s29[2],s28[2],s27[2],s26[2],s25[2],s24[2],s23[2],s22[2],s21[2],s20[2],s19[2],s18[2],s17[2],s16[2],s15[2],s14[2],s13[2],s12[2],s11[2],s10[2],s9[2],s8[2],s7[2],s6[2],s5[2],s4[2],s3[2],s2[2],s1[2],s0[2],ReadAd1,ReadData1[2]),
         m3 (s31[3],s30[3],s29[3],s28[3],s27[3],s26[3],s25[3],s24[3],s23[3],s22[3],s21[3],s20[3],s19[3],s18[3],s17[3],s16[3],s15[3],s14[3],s13[3],s12[3],s11[3],s10[3],s9[3],s8[3],s7[3],s6[3],s5[3],s4[3],s3[3],s2[3],s1[3],s0[3],ReadAd1,ReadData1[3]),
         m4 (s31[4],s30[4],s29[4],s28[4],s27[4],s26[4],s25[4],s24[4],s23[4],s22[4],s21[4],s20[4],s19[4],s18[4],s17[4],s16[4],s15[4],s14[4],s13[4],s12[4],s11[4],s10[4],s9[4],s8[4],s7[4],s6[4],s5[4],s4[4],s3[4],s2[4],s1[4],s0[4],ReadAd1,ReadData1[4]),
         m5 (s31[5],s30[5],s29[5],s28[5],s27[5],s26[5],s25[5],s24[5],s23[5],s22[5],s21[5],s20[5],s19[5],s18[5],s17[5],s16[5],s15[5],s14[5],s13[5],s12[5],s11[5],s10[5],s9[5],s8[5],s7[5],s6[5],s5[5],s4[5],s3[5],s2[5],s1[5],s0[5],ReadAd1,ReadData1[5]),
         m6 (s31[6],s30[6],s29[6],s28[6],s27[6],s26[6],s25[6],s24[6],s23[6],s22[6],s21[6],s20[6],s19[6],s18[6],s17[6],s16[6],s15[6],s14[6],s13[6],s12[6],s11[6],s10[6],s9[6],s8[6],s7[6],s6[6],s5[6],s4[6],s3[6],s2[6],s1[6],s0[6],ReadAd1,ReadData1[6]),
         m7 (s31[7],s30[7],s29[7],s28[7],s27[7],s26[7],s25[7],s24[7],s23[7],s22[7],s21[7],s20[7],s19[7],s18[7],s17[7],s16[7],s15[7],s14[7],s13[7],s12[7],s11[7],s10[7],s9[7],s8[7],s7[7],s6[7],s5[7],s4[7],s3[7],s2[7],s1[7],s0[7],ReadAd1,ReadData1[7]),
         m8 (s31[8],s30[8],s29[8],s28[8],s27[8],s26[8],s25[8],s24[8],s23[8],s22[8],s21[8],s20[8],s19[8],s18[8],s17[8],s16[8],s15[8],s14[8],s13[8],s12[8],s11[8],s10[8],s9[8],s8[8],s7[8],s6[8],s5[8],s4[8],s3[8],s2[8],s1[8],s0[8],ReadAd1,ReadData1[8]),
         m9 (s31[9],s30[9],s29[9],s28[9],s27[9],s26[9],s25[9],s24[9],s23[9],s22[9],s21[9],s20[9],s19[9],s18[9],s17[9],s16[9],s15[9],s14[9],s13[9],s12[9],s11[9],s10[9],s9[9],s8[9],s7[9],s6[9],s5[9],s4[9],s3[9],s2[9],s1[9],s0[9],ReadAd1,ReadData1[9]),
         m10 (s31[10],s30[10],s29[10],s28[10],s27[10],s26[10],s25[10],s24[10],s23[10],s22[10],s21[10],s20[10],s19[10],s18[10],s17[10],s16[10],s15[10],s14[10],s13[10],s12[10],s11[10],s10[10],s9[10],s8[10],s7[10],s6[10],s5[10],s4[10],s3[10],s2[10],s1[10],s0[10],ReadAd1,ReadData1[10]),
         m11 (s31[11],s30[11],s29[11],s28[11],s27[11],s26[11],s25[11],s24[11],s23[11],s22[11],s21[11],s20[11],s19[11],s18[11],s17[11],s16[11],s15[11],s14[11],s13[11],s12[11],s11[11],s10[11],s9[11],s8[11],s7[11],s6[11],s5[11],s4[11],s3[11],s2[11],s1[11],s0[11],ReadAd1,ReadData1[11]),
         m12 (s31[12],s30[12],s29[12],s28[12],s27[12],s26[12],s25[12],s24[12],s23[12],s22[12],s21[12],s20[12],s19[12],s18[12],s17[12],s16[12],s15[12],s14[12],s13[12],s12[12],s11[12],s10[12],s9[12],s8[12],s7[12],s6[12],s5[12],s4[12],s3[12],s2[12],s1[12],s0[12],ReadAd1,ReadData1[12]),
         m13 (s31[13],s30[13],s29[13],s28[13],s27[13],s26[13],s25[13],s24[13],s23[13],s22[13],s21[13],s20[13],s19[13],s18[13],s17[13],s16[13],s15[13],s14[13],s13[13],s12[13],s11[13],s10[13],s9[13],s8[13],s7[13],s6[13],s5[13],s4[13],s3[13],s2[13],s1[13],s0[13],ReadAd1,ReadData1[13]),
         m14 (s31[14],s30[14],s29[14],s28[14],s27[14],s26[14],s25[14],s24[14],s23[14],s22[14],s21[14],s20[14],s19[14],s18[14],s17[14],s16[14],s15[14],s14[14],s13[14],s12[14],s11[14],s10[14],s9[14],s8[14],s7[14],s6[14],s5[14],s4[14],s3[14],s2[14],s1[14],s0[14],ReadAd1,ReadData1[14]),
         m15 (s31[15],s30[15],s29[15],s28[15],s27[15],s26[15],s25[15],s24[15],s23[15],s22[15],s21[15],s20[15],s19[15],s18[15],s17[15],s16[15],s15[15],s14[15],s13[15],s12[15],s11[15],s10[15],s9[15],s8[15],s7[15],s6[15],s5[15],s4[15],s3[15],s2[15],s1[15],s0[15],ReadAd1,ReadData1[15]),
         m16 (s31[16],s30[16],s29[16],s28[16],s27[16],s26[16],s25[16],s24[16],s23[16],s22[16],s21[16],s20[16],s19[16],s18[16],s17[16],s16[16],s15[16],s14[16],s13[16],s12[16],s11[16],s10[16],s9[16],s8[16],s7[16],s6[16],s5[16],s4[16],s3[16],s2[16],s1[16],s0[16],ReadAd1,ReadData1[16]),
         m17 (s31[17],s30[17],s29[17],s28[17],s27[17],s26[17],s25[17],s24[17],s23[17],s22[17],s21[17],s20[17],s19[17],s18[17],s17[17],s16[17],s15[17],s14[17],s13[17],s12[17],s11[17],s10[17],s9[17],s8[17],s7[17],s6[17],s5[17],s4[17],s3[17],s2[17],s1[17],s0[17],ReadAd1,ReadData1[17]),
         m18 (s31[18],s30[18],s29[18],s28[18],s27[18],s26[18],s25[18],s24[18],s23[18],s22[18],s21[18],s20[18],s19[18],s18[18],s17[18],s16[18],s15[18],s14[18],s13[18],s12[18],s11[18],s10[18],s9[18],s8[18],s7[18],s6[18],s5[18],s4[18],s3[18],s2[18],s1[18],s0[18],ReadAd1,ReadData1[18]),
         m19 (s31[19],s30[19],s29[19],s28[19],s27[19],s26[19],s25[19],s24[19],s23[19],s22[19],s21[19],s20[19],s19[19],s18[19],s17[19],s16[19],s15[19],s14[19],s13[19],s12[19],s11[19],s10[19],s9[19],s8[19],s7[19],s6[19],s5[19],s4[19],s3[19],s2[19],s1[19],s0[19],ReadAd1,ReadData1[19]),
         m20 (s31[20],s30[20],s29[20],s28[20],s27[20],s26[20],s25[20],s24[20],s23[20],s22[20],s21[20],s20[20],s19[20],s18[20],s17[20],s16[20],s15[20],s14[20],s13[20],s12[20],s11[20],s10[20],s9[20],s8[20],s7[20],s6[20],s5[20],s4[20],s3[20],s2[20],s1[20],s0[20],ReadAd1,ReadData1[20]),
         m21 (s31[21],s30[21],s29[21],s28[21],s27[21],s26[21],s25[21],s24[21],s23[21],s22[21],s21[21],s20[21],s19[21],s18[21],s17[21],s16[21],s15[21],s14[21],s13[21],s12[21],s11[21],s10[21],s9[21],s8[21],s7[21],s6[21],s5[21],s4[21],s3[21],s2[21],s1[21],s0[21],ReadAd1,ReadData1[21]),
         m22 (s31[22],s30[22],s29[22],s28[22],s27[22],s26[22],s25[22],s24[22],s23[22],s22[22],s21[22],s20[22],s19[22],s18[22],s17[22],s16[22],s15[22],s14[22],s13[22],s12[22],s11[22],s10[22],s9[22],s8[22],s7[22],s6[22],s5[22],s4[22],s3[22],s2[22],s1[22],s0[22],ReadAd1,ReadData1[22]),
         m23 (s31[23],s30[23],s29[23],s28[23],s27[23],s26[23],s25[23],s24[23],s23[23],s22[23],s21[23],s20[23],s19[23],s18[23],s17[23],s16[23],s15[23],s14[23],s13[23],s12[23],s11[23],s10[23],s9[23],s8[23],s7[23],s6[23],s5[23],s4[23],s3[23],s2[23],s1[23],s0[23],ReadAd1,ReadData1[23]),
         m24 (s31[24],s30[24],s29[24],s28[24],s27[24],s26[24],s25[24],s24[24],s23[24],s22[24],s21[24],s20[24],s19[24],s18[24],s17[24],s16[24],s15[24],s14[24],s13[24],s12[24],s11[24],s10[24],s9[24],s8[24],s7[24],s6[24],s5[24],s4[24],s3[24],s2[24],s1[24],s0[24],ReadAd1,ReadData1[24]),
         m25 (s31[25],s30[25],s29[25],s28[25],s27[25],s26[25],s25[25],s24[25],s23[25],s22[25],s21[25],s20[25],s19[25],s18[25],s17[25],s16[25],s15[25],s14[25],s13[25],s12[25],s11[25],s10[25],s9[25],s8[25],s7[25],s6[25],s5[25],s4[25],s3[25],s2[25],s1[25],s0[25],ReadAd1,ReadData1[25]),
         m26 (s31[26],s30[26],s29[26],s28[26],s27[26],s26[26],s25[26],s24[26],s23[26],s22[26],s21[26],s20[26],s19[26],s18[26],s17[26],s16[26],s15[26],s14[26],s13[26],s12[26],s11[26],s10[26],s9[26],s8[26],s7[26],s6[26],s5[26],s4[26],s3[26],s2[26],s1[26],s0[26],ReadAd1,ReadData1[26]),
         m27 (s31[27],s30[27],s29[27],s28[27],s27[27],s26[27],s25[27],s24[27],s23[27],s22[27],s21[27],s20[27],s19[27],s18[27],s17[27],s16[27],s15[27],s14[27],s13[27],s12[27],s11[27],s10[27],s9[27],s8[27],s7[27],s6[27],s5[27],s4[27],s3[27],s2[27],s1[27],s0[27],ReadAd1,ReadData1[27]),
         m28 (s31[28],s30[28],s29[28],s28[28],s27[28],s26[28],s25[28],s24[28],s23[28],s22[28],s21[28],s20[28],s19[28],s18[28],s17[28],s16[28],s15[28],s14[28],s13[28],s12[28],s11[28],s10[28],s9[28],s8[28],s7[28],s6[28],s5[28],s4[28],s3[28],s2[28],s1[28],s0[28],ReadAd1,ReadData1[28]),
         m29 (s31[29],s30[29],s29[29],s28[29],s27[29],s26[29],s25[29],s24[29],s23[29],s22[29],s21[29],s20[29],s19[29],s18[29],s17[29],s16[29],s15[29],s14[29],s13[29],s12[29],s11[29],s10[29],s9[29],s8[29],s7[29],s6[29],s5[29],s4[29],s3[29],s2[29],s1[29],s0[29],ReadAd1,ReadData1[29]),
         m30 (s31[30],s30[30],s29[30],s28[30],s27[30],s26[30],s25[30],s24[30],s23[30],s22[30],s21[30],s20[30],s19[30],s18[30],s17[30],s16[30],s15[30],s14[30],s13[30],s12[30],s11[30],s10[30],s9[30],s8[30],s7[30],s6[30],s5[30],s4[30],s3[30],s2[30],s1[30],s0[30],ReadAd1,ReadData1[30]),
         m31 (s31[31],s30[31],s29[31],s28[31],s27[31],s26[31],s25[31],s24[31],s23[31],s22[31],s21[31],s20[31],s19[31],s18[31],s17[31],s16[31],s15[31],s14[31],s13[31],s12[31],s11[31],s10[31],s9[31],s8[31],s7[31],s6[31],s5[31],s4[31],s3[31],s2[31],s1[31],s0[31],ReadAd1,ReadData1[31]),
         n0 (s31[0],s30[0],s29[0],s28[0],s27[0],s26[0],s25[0],s24[0],s23[0],s22[0],s21[0],s20[0],s19[0],s18[0],s17[0],s16[0],s15[0],s14[0],s13[0],s12[0],s11[0],s10[0],s9[0],s8[0],s7[0],s6[0],s5[0],s4[0],s3[0],s2[0],s1[0],s0[0],ReadAd2,ReadData2[0]),
         n1 (s31[1],s30[1],s29[1],s28[1],s27[1],s26[1],s25[1],s24[1],s23[1],s22[1],s21[1],s20[1],s19[1],s18[1],s17[1],s16[1],s15[1],s14[1],s13[1],s12[1],s11[1],s10[1],s9[1],s8[1],s7[1],s6[1],s5[1],s4[1],s3[1],s2[1],s1[1],s0[1],ReadAd2,ReadData2[1]),
         n2 (s31[2],s30[2],s29[2],s28[2],s27[2],s26[2],s25[2],s24[2],s23[2],s22[2],s21[2],s20[2],s19[2],s18[2],s17[2],s16[2],s15[2],s14[2],s13[2],s12[2],s11[2],s10[2],s9[2],s8[2],s7[2],s6[2],s5[2],s4[2],s3[2],s2[2],s1[2],s0[2],ReadAd2,ReadData2[2]),
         n3 (s31[3],s30[3],s29[3],s28[3],s27[3],s26[3],s25[3],s24[3],s23[3],s22[3],s21[3],s20[3],s19[3],s18[3],s17[3],s16[3],s15[3],s14[3],s13[3],s12[3],s11[3],s10[3],s9[3],s8[3],s7[3],s6[3],s5[3],s4[3],s3[3],s2[3],s1[3],s0[3],ReadAd2,ReadData2[3]),
         n4 (s31[4],s30[4],s29[4],s28[4],s27[4],s26[4],s25[4],s24[4],s23[4],s22[4],s21[4],s20[4],s19[4],s18[4],s17[4],s16[4],s15[4],s14[4],s13[4],s12[4],s11[4],s10[4],s9[4],s8[4],s7[4],s6[4],s5[4],s4[4],s3[4],s2[4],s1[4],s0[4],ReadAd2,ReadData2[4]),
         n5 (s31[5],s30[5],s29[5],s28[5],s27[5],s26[5],s25[5],s24[5],s23[5],s22[5],s21[5],s20[5],s19[5],s18[5],s17[5],s16[5],s15[5],s14[5],s13[5],s12[5],s11[5],s10[5],s9[5],s8[5],s7[5],s6[5],s5[5],s4[5],s3[5],s2[5],s1[5],s0[5],ReadAd2,ReadData2[5]),
         n6 (s31[6],s30[6],s29[6],s28[6],s27[6],s26[6],s25[6],s24[6],s23[6],s22[6],s21[6],s20[6],s19[6],s18[6],s17[6],s16[6],s15[6],s14[6],s13[6],s12[6],s11[6],s10[6],s9[6],s8[6],s7[6],s6[6],s5[6],s4[6],s3[6],s2[6],s1[6],s0[6],ReadAd2,ReadData2[6]),
         n7 (s31[7],s30[7],s29[7],s28[7],s27[7],s26[7],s25[7],s24[7],s23[7],s22[7],s21[7],s20[7],s19[7],s18[7],s17[7],s16[7],s15[7],s14[7],s13[7],s12[7],s11[7],s10[7],s9[7],s8[7],s7[7],s6[7],s5[7],s4[7],s3[7],s2[7],s1[7],s0[7],ReadAd2,ReadData2[7]),
         n8 (s31[8],s30[8],s29[8],s28[8],s27[8],s26[8],s25[8],s24[8],s23[8],s22[8],s21[8],s20[8],s19[8],s18[8],s17[8],s16[8],s15[8],s14[8],s13[8],s12[8],s11[8],s10[8],s9[8],s8[8],s7[8],s6[8],s5[8],s4[8],s3[8],s2[8],s1[8],s0[8],ReadAd2,ReadData2[8]),
         n9 (s31[9],s30[9],s29[9],s28[9],s27[9],s26[9],s25[9],s24[9],s23[9],s22[9],s21[9],s20[9],s19[9],s18[9],s17[9],s16[9],s15[9],s14[9],s13[9],s12[9],s11[9],s10[9],s9[9],s8[9],s7[9],s6[9],s5[9],s4[9],s3[9],s2[9],s1[9],s0[9],ReadAd2,ReadData2[9]),
         n10 (s31[10],s30[10],s29[10],s28[10],s27[10],s26[10],s25[10],s24[10],s23[10],s22[10],s21[10],s20[10],s19[10],s18[10],s17[10],s16[10],s15[10],s14[10],s13[10],s12[10],s11[10],s10[10],s9[10],s8[10],s7[10],s6[10],s5[10],s4[10],s3[10],s2[10],s1[10],s0[10],ReadAd2,ReadData2[10]),
         n11 (s31[11],s30[11],s29[11],s28[11],s27[11],s26[11],s25[11],s24[11],s23[11],s22[11],s21[11],s20[11],s19[11],s18[11],s17[11],s16[11],s15[11],s14[11],s13[11],s12[11],s11[11],s10[11],s9[11],s8[11],s7[11],s6[11],s5[11],s4[11],s3[11],s2[11],s1[11],s0[11],ReadAd2,ReadData2[11]),
         n12 (s31[12],s30[12],s29[12],s28[12],s27[12],s26[12],s25[12],s24[12],s23[12],s22[12],s21[12],s20[12],s19[12],s18[12],s17[12],s16[12],s15[12],s14[12],s13[12],s12[12],s11[12],s10[12],s9[12],s8[12],s7[12],s6[12],s5[12],s4[12],s3[12],s2[12],s1[12],s0[12],ReadAd2,ReadData2[12]),
         n13 (s31[13],s30[13],s29[13],s28[13],s27[13],s26[13],s25[13],s24[13],s23[13],s22[13],s21[13],s20[13],s19[13],s18[13],s17[13],s16[13],s15[13],s14[13],s13[13],s12[13],s11[13],s10[13],s9[13],s8[13],s7[13],s6[13],s5[13],s4[13],s3[13],s2[13],s1[13],s0[13],ReadAd2,ReadData2[13]),
         n14 (s31[14],s30[14],s29[14],s28[14],s27[14],s26[14],s25[14],s24[14],s23[14],s22[14],s21[14],s20[14],s19[14],s18[14],s17[14],s16[14],s15[14],s14[14],s13[14],s12[14],s11[14],s10[14],s9[14],s8[14],s7[14],s6[14],s5[14],s4[14],s3[14],s2[14],s1[14],s0[14],ReadAd2,ReadData2[14]),
         n15 (s31[15],s30[15],s29[15],s28[15],s27[15],s26[15],s25[15],s24[15],s23[15],s22[15],s21[15],s20[15],s19[15],s18[15],s17[15],s16[15],s15[15],s14[15],s13[15],s12[15],s11[15],s10[15],s9[15],s8[15],s7[15],s6[15],s5[15],s4[15],s3[15],s2[15],s1[15],s0[15],ReadAd2,ReadData2[15]),
         n16 (s31[16],s30[16],s29[16],s28[16],s27[16],s26[16],s25[16],s24[16],s23[16],s22[16],s21[16],s20[16],s19[16],s18[16],s17[16],s16[16],s15[16],s14[16],s13[16],s12[16],s11[16],s10[16],s9[16],s8[16],s7[16],s6[16],s5[16],s4[16],s3[16],s2[16],s1[16],s0[16],ReadAd2,ReadData2[16]),
         n17 (s31[17],s30[17],s29[17],s28[17],s27[17],s26[17],s25[17],s24[17],s23[17],s22[17],s21[17],s20[17],s19[17],s18[17],s17[17],s16[17],s15[17],s14[17],s13[17],s12[17],s11[17],s10[17],s9[17],s8[17],s7[17],s6[17],s5[17],s4[17],s3[17],s2[17],s1[17],s0[17],ReadAd2,ReadData2[17]),
         n18 (s31[18],s30[18],s29[18],s28[18],s27[18],s26[18],s25[18],s24[18],s23[18],s22[18],s21[18],s20[18],s19[18],s18[18],s17[18],s16[18],s15[18],s14[18],s13[18],s12[18],s11[18],s10[18],s9[18],s8[18],s7[18],s6[18],s5[18],s4[18],s3[18],s2[18],s1[18],s0[18],ReadAd2,ReadData2[18]),
         n19 (s31[19],s30[19],s29[19],s28[19],s27[19],s26[19],s25[19],s24[19],s23[19],s22[19],s21[19],s20[19],s19[19],s18[19],s17[19],s16[19],s15[19],s14[19],s13[19],s12[19],s11[19],s10[19],s9[19],s8[19],s7[19],s6[19],s5[19],s4[19],s3[19],s2[19],s1[19],s0[19],ReadAd2,ReadData2[19]),
         n20 (s31[20],s30[20],s29[20],s28[20],s27[20],s26[20],s25[20],s24[20],s23[20],s22[20],s21[20],s20[20],s19[20],s18[20],s17[20],s16[20],s15[20],s14[20],s13[20],s12[20],s11[20],s10[20],s9[20],s8[20],s7[20],s6[20],s5[20],s4[20],s3[20],s2[20],s1[20],s0[20],ReadAd2,ReadData2[20]),
         n21 (s31[21],s30[21],s29[21],s28[21],s27[21],s26[21],s25[21],s24[21],s23[21],s22[21],s21[21],s20[21],s19[21],s18[21],s17[21],s16[21],s15[21],s14[21],s13[21],s12[21],s11[21],s10[21],s9[21],s8[21],s7[21],s6[21],s5[21],s4[21],s3[21],s2[21],s1[21],s0[21],ReadAd2,ReadData2[21]),
         n22 (s31[22],s30[22],s29[22],s28[22],s27[22],s26[22],s25[22],s24[22],s23[22],s22[22],s21[22],s20[22],s19[22],s18[22],s17[22],s16[22],s15[22],s14[22],s13[22],s12[22],s11[22],s10[22],s9[22],s8[22],s7[22],s6[22],s5[22],s4[22],s3[22],s2[22],s1[22],s0[22],ReadAd2,ReadData2[22]),
         n23 (s31[23],s30[23],s29[23],s28[23],s27[23],s26[23],s25[23],s24[23],s23[23],s22[23],s21[23],s20[23],s19[23],s18[23],s17[23],s16[23],s15[23],s14[23],s13[23],s12[23],s11[23],s10[23],s9[23],s8[23],s7[23],s6[23],s5[23],s4[23],s3[23],s2[23],s1[23],s0[23],ReadAd2,ReadData2[23]),
         n24 (s31[24],s30[24],s29[24],s28[24],s27[24],s26[24],s25[24],s24[24],s23[24],s22[24],s21[24],s20[24],s19[24],s18[24],s17[24],s16[24],s15[24],s14[24],s13[24],s12[24],s11[24],s10[24],s9[24],s8[24],s7[24],s6[24],s5[24],s4[24],s3[24],s2[24],s1[24],s0[24],ReadAd2,ReadData2[24]),
         n25 (s31[25],s30[25],s29[25],s28[25],s27[25],s26[25],s25[25],s24[25],s23[25],s22[25],s21[25],s20[25],s19[25],s18[25],s17[25],s16[25],s15[25],s14[25],s13[25],s12[25],s11[25],s10[25],s9[25],s8[25],s7[25],s6[25],s5[25],s4[25],s3[25],s2[25],s1[25],s0[25],ReadAd2,ReadData2[25]),
         n26 (s31[26],s30[26],s29[26],s28[26],s27[26],s26[26],s25[26],s24[26],s23[26],s22[26],s21[26],s20[26],s19[26],s18[26],s17[26],s16[26],s15[26],s14[26],s13[26],s12[26],s11[26],s10[26],s9[26],s8[26],s7[26],s6[26],s5[26],s4[26],s3[26],s2[26],s1[26],s0[26],ReadAd2,ReadData2[26]),
         n27 (s31[27],s30[27],s29[27],s28[27],s27[27],s26[27],s25[27],s24[27],s23[27],s22[27],s21[27],s20[27],s19[27],s18[27],s17[27],s16[27],s15[27],s14[27],s13[27],s12[27],s11[27],s10[27],s9[27],s8[27],s7[27],s6[27],s5[27],s4[27],s3[27],s2[27],s1[27],s0[27],ReadAd2,ReadData2[27]),
         n28 (s31[28],s30[28],s29[28],s28[28],s27[28],s26[28],s25[28],s24[28],s23[28],s22[28],s21[28],s20[28],s19[28],s18[28],s17[28],s16[28],s15[28],s14[28],s13[28],s12[28],s11[28],s10[28],s9[28],s8[28],s7[28],s6[28],s5[28],s4[28],s3[28],s2[28],s1[28],s0[28],ReadAd2,ReadData2[28]),
         n29 (s31[29],s30[29],s29[29],s28[29],s27[29],s26[29],s25[29],s24[29],s23[29],s22[29],s21[29],s20[29],s19[29],s18[29],s17[29],s16[29],s15[29],s14[29],s13[29],s12[29],s11[29],s10[29],s9[29],s8[29],s7[29],s6[29],s5[29],s4[29],s3[29],s2[29],s1[29],s0[29],ReadAd2,ReadData2[29]),
         n30 (s31[30],s30[30],s29[30],s28[30],s27[30],s26[30],s25[30],s24[30],s23[30],s22[30],s21[30],s20[30],s19[30],s18[30],s17[30],s16[30],s15[30],s14[30],s13[30],s12[30],s11[30],s10[30],s9[30],s8[30],s7[30],s6[30],s5[30],s4[30],s3[30],s2[30],s1[30],s0[30],ReadAd2,ReadData2[30]),
         n31 (s31[31],s30[31],s29[31],s28[31],s27[31],s26[31],s25[31],s24[31],s23[31],s22[31],s21[31],s20[31],s19[31],s18[31],s17[31],s16[31],s15[31],s14[31],s13[31],s12[31],s11[31],s10[31],s9[31],s8[31],s7[31],s6[31],s5[31],s4[31],s3[31],s2[31],s1[31],s0[31],ReadAd2,ReadData2[31]),
         p0 (s31[0],s30[0],s29[0],s28[0],s27[0],s26[0],s25[0],s24[0],s23[0],s22[0],s21[0],s20[0],s19[0],s18[0],s17[0],s16[0],s15[0],s14[0],s13[0],s12[0],s11[0],s10[0],s9[0],s8[0],s7[0],s6[0],s5[0],s4[0],s3[0],s2[0],s1[0],s0[0],5'b11111,ReadData3[0]),
         p1 (s31[1],s30[1],s29[1],s28[1],s27[1],s26[1],s25[1],s24[1],s23[1],s22[1],s21[1],s20[1],s19[1],s18[1],s17[1],s16[1],s15[1],s14[1],s13[1],s12[1],s11[1],s10[1],s9[1],s8[1],s7[1],s6[1],s5[1],s4[1],s3[1],s2[1],s1[1],s0[1],5'b11111,ReadData3[1]),
         p2 (s31[2],s30[2],s29[2],s28[2],s27[2],s26[2],s25[2],s24[2],s23[2],s22[2],s21[2],s20[2],s19[2],s18[2],s17[2],s16[2],s15[2],s14[2],s13[2],s12[2],s11[2],s10[2],s9[2],s8[2],s7[2],s6[2],s5[2],s4[2],s3[2],s2[2],s1[2],s0[2],5'b11111,ReadData3[2]),
         p3 (s31[3],s30[3],s29[3],s28[3],s27[3],s26[3],s25[3],s24[3],s23[3],s22[3],s21[3],s20[3],s19[3],s18[3],s17[3],s16[3],s15[3],s14[3],s13[3],s12[3],s11[3],s10[3],s9[3],s8[3],s7[3],s6[3],s5[3],s4[3],s3[3],s2[3],s1[3],s0[3],5'b11111,ReadData3[3]),
         p4 (s31[4],s30[4],s29[4],s28[4],s27[4],s26[4],s25[4],s24[4],s23[4],s22[4],s21[4],s20[4],s19[4],s18[4],s17[4],s16[4],s15[4],s14[4],s13[4],s12[4],s11[4],s10[4],s9[4],s8[4],s7[4],s6[4],s5[4],s4[4],s3[4],s2[4],s1[4],s0[4],5'b11111,ReadData3[4]),
         p5 (s31[5],s30[5],s29[5],s28[5],s27[5],s26[5],s25[5],s24[5],s23[5],s22[5],s21[5],s20[5],s19[5],s18[5],s17[5],s16[5],s15[5],s14[5],s13[5],s12[5],s11[5],s10[5],s9[5],s8[5],s7[5],s6[5],s5[5],s4[5],s3[5],s2[5],s1[5],s0[5],5'b11111,ReadData3[5]),
         p6 (s31[6],s30[6],s29[6],s28[6],s27[6],s26[6],s25[6],s24[6],s23[6],s22[6],s21[6],s20[6],s19[6],s18[6],s17[6],s16[6],s15[6],s14[6],s13[6],s12[6],s11[6],s10[6],s9[6],s8[6],s7[6],s6[6],s5[6],s4[6],s3[6],s2[6],s1[6],s0[6],5'b11111,ReadData3[6]),
         p7 (s31[7],s30[7],s29[7],s28[7],s27[7],s26[7],s25[7],s24[7],s23[7],s22[7],s21[7],s20[7],s19[7],s18[7],s17[7],s16[7],s15[7],s14[7],s13[7],s12[7],s11[7],s10[7],s9[7],s8[7],s7[7],s6[7],s5[7],s4[7],s3[7],s2[7],s1[7],s0[7],5'b11111,ReadData3[7]),
         p8 (s31[8],s30[8],s29[8],s28[8],s27[8],s26[8],s25[8],s24[8],s23[8],s22[8],s21[8],s20[8],s19[8],s18[8],s17[8],s16[8],s15[8],s14[8],s13[8],s12[8],s11[8],s10[8],s9[8],s8[8],s7[8],s6[8],s5[8],s4[8],s3[8],s2[8],s1[8],s0[8],5'b11111,ReadData3[8]),
         p9 (s31[9],s30[9],s29[9],s28[9],s27[9],s26[9],s25[9],s24[9],s23[9],s22[9],s21[9],s20[9],s19[9],s18[9],s17[9],s16[9],s15[9],s14[9],s13[9],s12[9],s11[9],s10[9],s9[9],s8[9],s7[9],s6[9],s5[9],s4[9],s3[9],s2[9],s1[9],s0[9],5'b11111,ReadData3[9]),
         p10 (s31[10],s30[10],s29[10],s28[10],s27[10],s26[10],s25[10],s24[10],s23[10],s22[10],s21[10],s20[10],s19[10],s18[10],s17[10],s16[10],s15[10],s14[10],s13[10],s12[10],s11[10],s10[10],s9[10],s8[10],s7[10],s6[10],s5[10],s4[10],s3[10],s2[10],s1[10],s0[10],5'b11111,ReadData3[10]),
         p11 (s31[11],s30[11],s29[11],s28[11],s27[11],s26[11],s25[11],s24[11],s23[11],s22[11],s21[11],s20[11],s19[11],s18[11],s17[11],s16[11],s15[11],s14[11],s13[11],s12[11],s11[11],s10[11],s9[11],s8[11],s7[11],s6[11],s5[11],s4[11],s3[11],s2[11],s1[11],s0[11],5'b11111,ReadData3[11]),
         p12 (s31[12],s30[12],s29[12],s28[12],s27[12],s26[12],s25[12],s24[12],s23[12],s22[12],s21[12],s20[12],s19[12],s18[12],s17[12],s16[12],s15[12],s14[12],s13[12],s12[12],s11[12],s10[12],s9[12],s8[12],s7[12],s6[12],s5[12],s4[12],s3[12],s2[12],s1[12],s0[12],5'b11111,ReadData3[12]),
         p13 (s31[13],s30[13],s29[13],s28[13],s27[13],s26[13],s25[13],s24[13],s23[13],s22[13],s21[13],s20[13],s19[13],s18[13],s17[13],s16[13],s15[13],s14[13],s13[13],s12[13],s11[13],s10[13],s9[13],s8[13],s7[13],s6[13],s5[13],s4[13],s3[13],s2[13],s1[13],s0[13],5'b11111,ReadData3[13]),
         p14 (s31[14],s30[14],s29[14],s28[14],s27[14],s26[14],s25[14],s24[14],s23[14],s22[14],s21[14],s20[14],s19[14],s18[14],s17[14],s16[14],s15[14],s14[14],s13[14],s12[14],s11[14],s10[14],s9[14],s8[14],s7[14],s6[14],s5[14],s4[14],s3[14],s2[14],s1[14],s0[14],5'b11111,ReadData3[14]),
         p15 (s31[15],s30[15],s29[15],s28[15],s27[15],s26[15],s25[15],s24[15],s23[15],s22[15],s21[15],s20[15],s19[15],s18[15],s17[15],s16[15],s15[15],s14[15],s13[15],s12[15],s11[15],s10[15],s9[15],s8[15],s7[15],s6[15],s5[15],s4[15],s3[15],s2[15],s1[15],s0[15],5'b11111,ReadData3[15]),
         p16 (s31[16],s30[16],s29[16],s28[16],s27[16],s26[16],s25[16],s24[16],s23[16],s22[16],s21[16],s20[16],s19[16],s18[16],s17[16],s16[16],s15[16],s14[16],s13[16],s12[16],s11[16],s10[16],s9[16],s8[16],s7[16],s6[16],s5[16],s4[16],s3[16],s2[16],s1[16],s0[16],5'b11111,ReadData3[16]),
         p17 (s31[17],s30[17],s29[17],s28[17],s27[17],s26[17],s25[17],s24[17],s23[17],s22[17],s21[17],s20[17],s19[17],s18[17],s17[17],s16[17],s15[17],s14[17],s13[17],s12[17],s11[17],s10[17],s9[17],s8[17],s7[17],s6[17],s5[17],s4[17],s3[17],s2[17],s1[17],s0[17],5'b11111,ReadData3[17]),
         p18 (s31[18],s30[18],s29[18],s28[18],s27[18],s26[18],s25[18],s24[18],s23[18],s22[18],s21[18],s20[18],s19[18],s18[18],s17[18],s16[18],s15[18],s14[18],s13[18],s12[18],s11[18],s10[18],s9[18],s8[18],s7[18],s6[18],s5[18],s4[18],s3[18],s2[18],s1[18],s0[18],5'b11111,ReadData3[18]),
         p19 (s31[19],s30[19],s29[19],s28[19],s27[19],s26[19],s25[19],s24[19],s23[19],s22[19],s21[19],s20[19],s19[19],s18[19],s17[19],s16[19],s15[19],s14[19],s13[19],s12[19],s11[19],s10[19],s9[19],s8[19],s7[19],s6[19],s5[19],s4[19],s3[19],s2[19],s1[19],s0[19],5'b11111,ReadData3[19]),
         p20 (s31[20],s30[20],s29[20],s28[20],s27[20],s26[20],s25[20],s24[20],s23[20],s22[20],s21[20],s20[20],s19[20],s18[20],s17[20],s16[20],s15[20],s14[20],s13[20],s12[20],s11[20],s10[20],s9[20],s8[20],s7[20],s6[20],s5[20],s4[20],s3[20],s2[20],s1[20],s0[20],5'b11111,ReadData3[20]),
         p21 (s31[21],s30[21],s29[21],s28[21],s27[21],s26[21],s25[21],s24[21],s23[21],s22[21],s21[21],s20[21],s19[21],s18[21],s17[21],s16[21],s15[21],s14[21],s13[21],s12[21],s11[21],s10[21],s9[21],s8[21],s7[21],s6[21],s5[21],s4[21],s3[21],s2[21],s1[21],s0[21],5'b11111,ReadData3[21]),
         p22 (s31[22],s30[22],s29[22],s28[22],s27[22],s26[22],s25[22],s24[22],s23[22],s22[22],s21[22],s20[22],s19[22],s18[22],s17[22],s16[22],s15[22],s14[22],s13[22],s12[22],s11[22],s10[22],s9[22],s8[22],s7[22],s6[22],s5[22],s4[22],s3[22],s2[22],s1[22],s0[22],5'b11111,ReadData3[22]),
         p23 (s31[23],s30[23],s29[23],s28[23],s27[23],s26[23],s25[23],s24[23],s23[23],s22[23],s21[23],s20[23],s19[23],s18[23],s17[23],s16[23],s15[23],s14[23],s13[23],s12[23],s11[23],s10[23],s9[23],s8[23],s7[23],s6[23],s5[23],s4[23],s3[23],s2[23],s1[23],s0[23],5'b11111,ReadData3[23]),
         p24 (s31[24],s30[24],s29[24],s28[24],s27[24],s26[24],s25[24],s24[24],s23[24],s22[24],s21[24],s20[24],s19[24],s18[24],s17[24],s16[24],s15[24],s14[24],s13[24],s12[24],s11[24],s10[24],s9[24],s8[24],s7[24],s6[24],s5[24],s4[24],s3[24],s2[24],s1[24],s0[24],5'b11111,ReadData3[24]),
         p25 (s31[25],s30[25],s29[25],s28[25],s27[25],s26[25],s25[25],s24[25],s23[25],s22[25],s21[25],s20[25],s19[25],s18[25],s17[25],s16[25],s15[25],s14[25],s13[25],s12[25],s11[25],s10[25],s9[25],s8[25],s7[25],s6[25],s5[25],s4[25],s3[25],s2[25],s1[25],s0[25],5'b11111,ReadData3[25]),
         p26 (s31[26],s30[26],s29[26],s28[26],s27[26],s26[26],s25[26],s24[26],s23[26],s22[26],s21[26],s20[26],s19[26],s18[26],s17[26],s16[26],s15[26],s14[26],s13[26],s12[26],s11[26],s10[26],s9[26],s8[26],s7[26],s6[26],s5[26],s4[26],s3[26],s2[26],s1[26],s0[26],5'b11111,ReadData3[26]),
         p27 (s31[27],s30[27],s29[27],s28[27],s27[27],s26[27],s25[27],s24[27],s23[27],s22[27],s21[27],s20[27],s19[27],s18[27],s17[27],s16[27],s15[27],s14[27],s13[27],s12[27],s11[27],s10[27],s9[27],s8[27],s7[27],s6[27],s5[27],s4[27],s3[27],s2[27],s1[27],s0[27],5'b11111,ReadData3[27]),
         p28 (s31[28],s30[28],s29[28],s28[28],s27[28],s26[28],s25[28],s24[28],s23[28],s22[28],s21[28],s20[28],s19[28],s18[28],s17[28],s16[28],s15[28],s14[28],s13[28],s12[28],s11[28],s10[28],s9[28],s8[28],s7[28],s6[28],s5[28],s4[28],s3[28],s2[28],s1[28],s0[28],5'b11111,ReadData3[28]),
         p29 (s31[29],s30[29],s29[29],s28[29],s27[29],s26[29],s25[29],s24[29],s23[29],s22[29],s21[29],s20[29],s19[29],s18[29],s17[29],s16[29],s15[29],s14[29],s13[29],s12[29],s11[29],s10[29],s9[29],s8[29],s7[29],s6[29],s5[29],s4[29],s3[29],s2[29],s1[29],s0[29],5'b11111,ReadData3[29]),
         p30 (s31[30],s30[30],s29[30],s28[30],s27[30],s26[30],s25[30],s24[30],s23[30],s22[30],s21[30],s20[30],s19[30],s18[30],s17[30],s16[30],s15[30],s14[30],s13[30],s12[30],s11[30],s10[30],s9[30],s8[30],s7[30],s6[30],s5[30],s4[30],s3[30],s2[30],s1[30],s0[30],5'b11111,ReadData3[30]),
         p31 (s31[31],s30[31],s29[31],s28[31],s27[31],s26[31],s25[31],s24[31],s23[31],s22[31],s21[31],s20[31],s19[31],s18[31],s17[31],s16[31],s15[31],s14[31],s13[31],s12[31],s11[31],s10[31],s9[31],s8[31],s7[31],s6[31],s5[31],s4[31],s3[31],s2[31],s1[31],s0[31],5'b11111,ReadData3[31]);
endmodule